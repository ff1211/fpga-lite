//****************************************************************
// Copyright 2023 Tianjin University 305 Lab. All Rights Reserved.
//
// File:
// control.sv
// 
// Description:
// Control module of remap core.
// 
// Revision history:
// Version  Date        Author      Changes      
// 1.0      2023.02.24  ff          Initial version
//****************************************************************

`timescale 1ns/1ps

module control #(
    parameter DATA_WIDTH = 16
) (
    input  logic    clk,
    input  logic    rst_n

);


    
endmodule